///////////////////////////////////////////////////
// HA.sv  This design will take in 2 bits       //
// and add them to produce a sum and carry     //
////////////////////////////////////////////////
module HA(
  input 	A,Cin,	// two input bits to be added
  output	S,Cout	// Sum and carry
);

	/////////////////////////////////////////////////
	// Declare any internal signals as type logic //
	///////////////////////////////////////////////
	
	/////////////////////////////////////////////////
	// Implement Half Adder as structural verilog //
	///////////////////////////////////////////////
	xor iXOR1(S,A,Cin);
	and iAND1(Cout,A,Cin);

endmodule